VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM256
  CLASS BLOCK ;
  FOREIGN RAM256 ;
  ORIGIN 0.000 0.000 ;
  SIZE 809.600 BY 533.120 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 807.600 55.800 809.600 56.400 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 807.600 93.880 809.600 94.480 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 807.600 131.960 809.600 132.560 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 807.600 170.040 809.600 170.640 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 807.600 208.120 809.600 208.720 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 807.600 246.200 809.600 246.800 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 807.600 284.280 809.600 284.880 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 807.600 322.360 809.600 322.960 ;
    END
  END A0[7]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 807.600 360.440 809.600 361.040 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 0.000 366.990 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 0.000 417.590 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 0.000 442.890 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 0.000 468.190 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 0.000 493.490 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 0.000 544.090 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.110 0.000 569.390 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 0.000 594.690 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 0.000 619.990 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 0.000 645.290 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 0.000 670.590 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.910 0.000 721.190 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 0.000 746.490 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 0.000 771.790 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.810 0.000 797.090 2.000 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 2.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 2.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 2.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 531.120 12.790 533.120 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 531.120 265.790 533.120 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 531.120 291.090 533.120 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 531.120 316.390 533.120 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 531.120 341.690 533.120 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 531.120 366.990 533.120 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 531.120 392.290 533.120 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 531.120 417.590 533.120 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 531.120 442.890 533.120 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 531.120 468.190 533.120 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 531.120 493.490 533.120 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 531.120 38.090 533.120 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 531.120 518.790 533.120 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 531.120 544.090 533.120 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.110 531.120 569.390 533.120 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 531.120 594.690 533.120 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 531.120 619.990 533.120 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 531.120 645.290 533.120 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 531.120 670.590 533.120 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 531.120 695.890 533.120 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.910 531.120 721.190 533.120 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 531.120 746.490 533.120 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 531.120 63.390 533.120 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 531.120 771.790 533.120 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.810 531.120 797.090 533.120 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 531.120 88.690 533.120 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 531.120 113.990 533.120 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 531.120 139.290 533.120 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 531.120 164.590 533.120 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 531.120 189.890 533.120 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 531.120 215.190 533.120 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 531.120 240.490 533.120 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 807.600 17.720 809.600 18.320 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 530.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.680 2.480 250.280 530.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 402.280 2.480 403.880 530.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 555.880 2.480 557.480 530.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 709.480 2.480 711.080 530.640 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 530.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 530.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 530.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 479.080 2.480 480.680 530.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.680 2.480 634.280 530.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.280 2.480 787.880 530.640 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 807.600 398.520 809.600 399.120 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 807.600 436.600 809.600 437.200 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 807.600 474.680 809.600 475.280 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 807.600 512.760 809.600 513.360 ;
    END
  END WE0[3]
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 806.840 530.485 ;
      LAYER met1 ;
        RECT 1.910 0.040 808.610 532.400 ;
      LAYER met2 ;
        RECT 1.010 530.840 12.230 532.965 ;
        RECT 13.070 530.840 37.530 532.965 ;
        RECT 38.370 530.840 62.830 532.965 ;
        RECT 63.670 530.840 88.130 532.965 ;
        RECT 88.970 530.840 113.430 532.965 ;
        RECT 114.270 530.840 138.730 532.965 ;
        RECT 139.570 530.840 164.030 532.965 ;
        RECT 164.870 530.840 189.330 532.965 ;
        RECT 190.170 530.840 214.630 532.965 ;
        RECT 215.470 530.840 239.930 532.965 ;
        RECT 240.770 530.840 265.230 532.965 ;
        RECT 266.070 530.840 290.530 532.965 ;
        RECT 291.370 530.840 315.830 532.965 ;
        RECT 316.670 530.840 341.130 532.965 ;
        RECT 341.970 530.840 366.430 532.965 ;
        RECT 367.270 530.840 391.730 532.965 ;
        RECT 392.570 530.840 417.030 532.965 ;
        RECT 417.870 530.840 442.330 532.965 ;
        RECT 443.170 530.840 467.630 532.965 ;
        RECT 468.470 530.840 492.930 532.965 ;
        RECT 493.770 530.840 518.230 532.965 ;
        RECT 519.070 530.840 543.530 532.965 ;
        RECT 544.370 530.840 568.830 532.965 ;
        RECT 569.670 530.840 594.130 532.965 ;
        RECT 594.970 530.840 619.430 532.965 ;
        RECT 620.270 530.840 644.730 532.965 ;
        RECT 645.570 530.840 670.030 532.965 ;
        RECT 670.870 530.840 695.330 532.965 ;
        RECT 696.170 530.840 720.630 532.965 ;
        RECT 721.470 530.840 745.930 532.965 ;
        RECT 746.770 530.840 771.230 532.965 ;
        RECT 772.070 530.840 796.530 532.965 ;
        RECT 797.370 530.840 808.580 532.965 ;
        RECT 1.010 2.280 808.580 530.840 ;
        RECT 1.010 0.010 12.230 2.280 ;
        RECT 13.070 0.010 37.530 2.280 ;
        RECT 38.370 0.010 62.830 2.280 ;
        RECT 63.670 0.010 88.130 2.280 ;
        RECT 88.970 0.010 113.430 2.280 ;
        RECT 114.270 0.010 138.730 2.280 ;
        RECT 139.570 0.010 164.030 2.280 ;
        RECT 164.870 0.010 189.330 2.280 ;
        RECT 190.170 0.010 214.630 2.280 ;
        RECT 215.470 0.010 239.930 2.280 ;
        RECT 240.770 0.010 265.230 2.280 ;
        RECT 266.070 0.010 290.530 2.280 ;
        RECT 291.370 0.010 315.830 2.280 ;
        RECT 316.670 0.010 341.130 2.280 ;
        RECT 341.970 0.010 366.430 2.280 ;
        RECT 367.270 0.010 391.730 2.280 ;
        RECT 392.570 0.010 417.030 2.280 ;
        RECT 417.870 0.010 442.330 2.280 ;
        RECT 443.170 0.010 467.630 2.280 ;
        RECT 468.470 0.010 492.930 2.280 ;
        RECT 493.770 0.010 518.230 2.280 ;
        RECT 519.070 0.010 543.530 2.280 ;
        RECT 544.370 0.010 568.830 2.280 ;
        RECT 569.670 0.010 594.130 2.280 ;
        RECT 594.970 0.010 619.430 2.280 ;
        RECT 620.270 0.010 644.730 2.280 ;
        RECT 645.570 0.010 670.030 2.280 ;
        RECT 670.870 0.010 695.330 2.280 ;
        RECT 696.170 0.010 720.630 2.280 ;
        RECT 721.470 0.010 745.930 2.280 ;
        RECT 746.770 0.010 771.230 2.280 ;
        RECT 772.070 0.010 796.530 2.280 ;
        RECT 797.370 0.010 808.580 2.280 ;
      LAYER met3 ;
        RECT 0.985 513.760 807.600 532.945 ;
        RECT 0.985 512.360 807.200 513.760 ;
        RECT 0.985 475.680 807.600 512.360 ;
        RECT 0.985 474.280 807.200 475.680 ;
        RECT 0.985 437.600 807.600 474.280 ;
        RECT 0.985 436.200 807.200 437.600 ;
        RECT 0.985 399.520 807.600 436.200 ;
        RECT 0.985 398.120 807.200 399.520 ;
        RECT 0.985 361.440 807.600 398.120 ;
        RECT 0.985 360.040 807.200 361.440 ;
        RECT 0.985 323.360 807.600 360.040 ;
        RECT 0.985 321.960 807.200 323.360 ;
        RECT 0.985 285.280 807.600 321.960 ;
        RECT 0.985 283.880 807.200 285.280 ;
        RECT 0.985 247.200 807.600 283.880 ;
        RECT 0.985 245.800 807.200 247.200 ;
        RECT 0.985 209.120 807.600 245.800 ;
        RECT 0.985 207.720 807.200 209.120 ;
        RECT 0.985 171.040 807.600 207.720 ;
        RECT 0.985 169.640 807.200 171.040 ;
        RECT 0.985 132.960 807.600 169.640 ;
        RECT 0.985 131.560 807.200 132.960 ;
        RECT 0.985 94.880 807.600 131.560 ;
        RECT 0.985 93.480 807.200 94.880 ;
        RECT 0.985 56.800 807.600 93.480 ;
        RECT 0.985 55.400 807.200 56.800 ;
        RECT 0.985 18.720 807.600 55.400 ;
        RECT 0.985 17.320 807.200 18.720 ;
        RECT 0.985 0.175 807.600 17.320 ;
      LAYER met4 ;
        RECT 38.935 5.615 94.680 526.825 ;
        RECT 97.080 5.615 171.480 526.825 ;
        RECT 173.880 5.615 248.280 526.825 ;
        RECT 250.680 5.615 325.080 526.825 ;
        RECT 327.480 5.615 401.880 526.825 ;
        RECT 404.280 5.615 478.680 526.825 ;
        RECT 481.080 5.615 555.480 526.825 ;
        RECT 557.880 5.615 632.280 526.825 ;
        RECT 634.680 5.615 709.080 526.825 ;
        RECT 711.480 5.615 785.880 526.825 ;
        RECT 788.280 5.615 800.105 526.825 ;
  END
END RAM256
END LIBRARY

