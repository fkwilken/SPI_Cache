VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM256
  CLASS BLOCK ;
  FOREIGN RAM256 ;
  ORIGIN 0.000 0.000 ;
  SIZE 434.240 BY 446.080 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 432.240 57.160 434.240 57.760 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 432.240 93.880 434.240 94.480 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 432.240 130.600 434.240 131.200 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 432.240 167.320 434.240 167.920 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 432.240 204.040 434.240 204.640 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 432.240 240.760 434.240 241.360 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 432.240 277.480 434.240 278.080 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 432.240 314.200 434.240 314.800 ;
    END
  END A0[7]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 432.240 350.920 434.240 351.520 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 2.000 ;
    END
  END Di0[15]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 2.000 ;
    END
  END Di0[1]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 2.000 ;
    END
  END Di0[2]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 2.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 2.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 2.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 444.080 13.710 446.080 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 444.080 285.110 446.080 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 444.080 312.250 446.080 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 444.080 339.390 446.080 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 444.080 366.530 446.080 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 444.080 393.670 446.080 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 444.080 420.810 446.080 ;
    END
  END Do0[15]
  PIN Do0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 444.080 40.850 446.080 ;
    END
  END Do0[1]
  PIN Do0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 444.080 67.990 446.080 ;
    END
  END Do0[2]
  PIN Do0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 444.080 95.130 446.080 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 444.080 122.270 446.080 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 444.080 149.410 446.080 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 444.080 176.550 446.080 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 444.080 203.690 446.080 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 444.080 230.830 446.080 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 444.080 257.970 446.080 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 432.240 20.440 434.240 21.040 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 443.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.680 2.480 250.280 443.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 402.280 2.480 403.880 443.600 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 443.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 443.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 443.600 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 432.240 387.640 434.240 388.240 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 432.240 424.360 434.240 424.960 ;
    END
  END WE0[1]
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 431.480 443.445 ;
      LAYER met1 ;
        RECT 2.370 0.720 433.250 446.040 ;
      LAYER met2 ;
        RECT 2.400 443.800 13.150 446.070 ;
        RECT 13.990 443.800 40.290 446.070 ;
        RECT 41.130 443.800 67.430 446.070 ;
        RECT 68.270 443.800 94.570 446.070 ;
        RECT 95.410 443.800 121.710 446.070 ;
        RECT 122.550 443.800 148.850 446.070 ;
        RECT 149.690 443.800 175.990 446.070 ;
        RECT 176.830 443.800 203.130 446.070 ;
        RECT 203.970 443.800 230.270 446.070 ;
        RECT 231.110 443.800 257.410 446.070 ;
        RECT 258.250 443.800 284.550 446.070 ;
        RECT 285.390 443.800 311.690 446.070 ;
        RECT 312.530 443.800 338.830 446.070 ;
        RECT 339.670 443.800 365.970 446.070 ;
        RECT 366.810 443.800 393.110 446.070 ;
        RECT 393.950 443.800 420.250 446.070 ;
        RECT 421.090 443.800 433.220 446.070 ;
        RECT 2.400 2.280 433.220 443.800 ;
        RECT 2.400 0.155 13.150 2.280 ;
        RECT 13.990 0.155 40.290 2.280 ;
        RECT 41.130 0.155 67.430 2.280 ;
        RECT 68.270 0.155 94.570 2.280 ;
        RECT 95.410 0.155 121.710 2.280 ;
        RECT 122.550 0.155 148.850 2.280 ;
        RECT 149.690 0.155 175.990 2.280 ;
        RECT 176.830 0.155 203.130 2.280 ;
        RECT 203.970 0.155 230.270 2.280 ;
        RECT 231.110 0.155 257.410 2.280 ;
        RECT 258.250 0.155 284.550 2.280 ;
        RECT 285.390 0.155 311.690 2.280 ;
        RECT 312.530 0.155 338.830 2.280 ;
        RECT 339.670 0.155 365.970 2.280 ;
        RECT 366.810 0.155 393.110 2.280 ;
        RECT 393.950 0.155 420.250 2.280 ;
        RECT 421.090 0.155 433.220 2.280 ;
      LAYER met3 ;
        RECT 2.825 425.360 432.240 443.525 ;
        RECT 2.825 423.960 431.840 425.360 ;
        RECT 2.825 388.640 432.240 423.960 ;
        RECT 2.825 387.240 431.840 388.640 ;
        RECT 2.825 351.920 432.240 387.240 ;
        RECT 2.825 350.520 431.840 351.920 ;
        RECT 2.825 315.200 432.240 350.520 ;
        RECT 2.825 313.800 431.840 315.200 ;
        RECT 2.825 278.480 432.240 313.800 ;
        RECT 2.825 277.080 431.840 278.480 ;
        RECT 2.825 241.760 432.240 277.080 ;
        RECT 2.825 240.360 431.840 241.760 ;
        RECT 2.825 205.040 432.240 240.360 ;
        RECT 2.825 203.640 431.840 205.040 ;
        RECT 2.825 168.320 432.240 203.640 ;
        RECT 2.825 166.920 431.840 168.320 ;
        RECT 2.825 131.600 432.240 166.920 ;
        RECT 2.825 130.200 431.840 131.600 ;
        RECT 2.825 94.880 432.240 130.200 ;
        RECT 2.825 93.480 431.840 94.880 ;
        RECT 2.825 58.160 432.240 93.480 ;
        RECT 2.825 56.760 431.840 58.160 ;
        RECT 2.825 21.440 432.240 56.760 ;
        RECT 2.825 20.040 431.840 21.440 ;
        RECT 2.825 0.175 432.240 20.040 ;
      LAYER met4 ;
        RECT 26.975 4.255 94.680 441.825 ;
        RECT 97.080 4.255 171.480 441.825 ;
        RECT 173.880 4.255 248.280 441.825 ;
        RECT 250.680 4.255 325.080 441.825 ;
        RECT 327.480 4.255 401.880 441.825 ;
        RECT 404.280 4.255 420.145 441.825 ;
  END
END RAM256
END LIBRARY

